entity b is
end b;

architecture struct of b is
begin
  a_inst: entity work.a;
end struct;
