entity old is
end old;
architecture behav of old is
begin
end behav;
