entity c is
end c;
architecture behav of c is
begin
end behav;
