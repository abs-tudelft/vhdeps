entity a is
end a;

architecture struct of a is
begin
  b_inst: entity work.b;
end struct;
