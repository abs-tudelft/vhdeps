-- Copyright 2018 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.TestCase_pkg.all;
use work.StreamSource_pkg.all;
use work.StreamSink_pkg.all;
use work.UtilInt_pkg.all;

entity StreamGearbox_tv is
end StreamGearbox_tv;

architecture TestVector of StreamGearbox_tv is
begin

  random_tc: process is
    constant TEST_STR : string(1 to 44) := "The quick brown fox jumps over the lazy dog.";
    variable a        : streamsource_type;
    variable b        : streamsink_type;
    variable remain   : integer;
    variable expect   : integer;
  begin
    tc_open("StreamGearbox-random",
      "tests that the data passes through unchanged with randomized timing and shape.");
    a.initialize("a");
    b.initialize("b");

    a.set_total_cyc(-5, 5);
    a.set_count(1, 2*a.g_count_max);
    a.set_last_greed(true);
    for i in 0 to 15 loop
      a.push_str(TEST_STR(1 to 44 - i));
      a.transmit;
    end loop;

    b.set_total_cyc(-5, 5);
    b.unblock;

    tc_wait_for(50 us);

    -- Check packet data.
    for i in 0 to 15 loop
      tc_check(b.pq_get_str, TEST_STR(1 to 44 - i));
    end loop;
    tc_check(b.pq_ready, false);

    tc_pass;
    wait;
  end process;

end TestVector;

