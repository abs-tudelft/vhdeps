entity a is
end a;
architecture behav of a is
begin
end behav;
