entity synthesis is
end synthesis;
architecture behav of synthesis is
begin
end behav;
