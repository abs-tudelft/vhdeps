package test_pkg is
  component test is
    generic (
      test: boolean := false;
    );
  end component;
end package;
