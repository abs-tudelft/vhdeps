entity test is
end test;
architecture behav of test is
begin
end behav;
