entity a is
end a;

architecture struct of a is
begin
end struct;

entity b is
end b;

architecture struct of b is
begin
end struct;
