entity b is
end b;
architecture behav of b is
begin
end behav;
