entity new is
end new;
architecture behav of new is
begin
end behav;
