entity synth_only is
end synth_only;

architecture struct of synth_only is
begin
end struct;
