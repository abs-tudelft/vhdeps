entity simulation is
end simulation;
architecture behav of simulation is
begin
end behav;
