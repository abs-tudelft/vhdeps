package test_pk is
  component test is
    generic (
      test: boolean := false;
    );
  end component;
end package;
