entity test is
  generic (
    test: boolean := false;
  );
end test;

architecture behav of test is
begin
end behav;
