entity test is
end test;

architecture struct of test is
begin
  synth_only_inst: entity work.synth_only;
end struct;
