entity b is
end b;

architecture struct of b is
begin
end struct;
